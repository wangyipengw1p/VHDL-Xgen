--------------------------------------------------
-- Creat time: 2019-05-31 22:55:50
-- Platform: Linux
-- Engineer: wangyipeng
-- University
-- Version
--------------------------------------------------



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;

entity t5 is
port(
	clk	: in	std_logic;
	rst	: in	std_logic;
	t2_t4	: in	std_logic_vector(7 downto 0);
	t5_o	: in	std_logic;
);
end entity;

architecture behaviral of t5 is

begin

end architecture;