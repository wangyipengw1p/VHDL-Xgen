--------------------------------------------------
-- Creat time: 2019-05-31 22:46:38
-- Platform: Linux
-- Engineer: wangyipeng
-- University
-- Version
--------------------------------------------------



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;
package testVXGen_pkg is 

end package;

package body testVXGen_pkg is

end package body;
